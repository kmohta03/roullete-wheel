module mipstoArduino (input [5:0], output [5:0]);
